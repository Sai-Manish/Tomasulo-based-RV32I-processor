// Top Module will have all the module integrated.